module tmds_8_to_10_bit(
	input wire [7:0] bits_in,
	input wire [9:0] bits_out
)

endmodule

module main(
	input wire clk,
	
	output wire led5,
	output wire led6
);
endmodule