module main(
	input wire clk,
	
	output wire led5,
	output wire led6
);
endmodule